module main

fn output_d2(deps []DependencyGraph) ![]string {
	return []string{}
}
